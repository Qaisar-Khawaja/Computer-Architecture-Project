// ----  Probes  ----
`define PROBE_ADDR assign_memory_addr_i
`define PROBE_DATA_IN   assign_memory_data_i
`define PROBE_DATA_OUT assign_memory_data_o
`define PROBE_READ_EN   assign_memory_read_en_i
`define PROBE_WRITE_EN  assign_memory_write_en_i

`define PROBE_F_PC assign_fetch_pc_o
`define PROBE_F_INSN assign_fetch_insn_o
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd1
// ----  Top module  ----
