// ----  Probes  ----
`define PROBE_F_PC    assign_f_pc
`define PROBE_F_INSN  assign_f_insn
`define PROBE_D_PC     assign_d_pc
`define PROBE_D_OPCODE assign_d_opcode
`define PROBE_D_RD     assign_d_rd
`define PROBE_D_FUNCT3 assign_d_funct3
`define PROBE_D_RS1    assign_d_rs1
`define PROBE_D_RS2    assign_d_rs2
`define PROBE_D_FUNCT7 assign_d_funct7
`define PROBE_D_IMM    assign_d_imm
`define PROBE_D_SHAMT  assign_d_shamt
`define PROBE_I_IMM    assign_i_imm
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd2
// ----  Top module  ----